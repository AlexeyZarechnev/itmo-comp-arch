module ternary_min(a, b, out);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule

module ternary_max(a, b, out);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule

module ternary_any(a, b, out);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule

module ternary_consensus(a, b, out);
  input [1:0] a
  input [1:0] b;
  output [1:0] out;
  // TODO: implementation
endmodule
